`include "flit.sv"

module vc_allocator#(
    parameter int LANES_PER_CHANNEL = 2,
    parameter int VC_DEPTH = 8
) (
)

endmodule
