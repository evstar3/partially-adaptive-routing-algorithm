`include "flit.sv"

module vc_allocator#(
    parameter int LANES_PER_CHANNEL = 2,
    parameter int VC_DEPTH = 5,
    parameter int FLIT_SIZE = 32
) (

)

endmodule
